module delay4 (
    input  wire clk,
    input  wire reset,   // ͬ����λ
    input  wire in,
    input  wire data,
    output reg  out
);

    reg [2:0] cnt;        // �� (in & data) ����Ϊ 1 �� clk ��
    reg [1:0] pulse_cnt;  // out �����ȼ�����2 clk��
    reg fired;             // �Ƿ��Ѿ���������������

    always @(posedge clk) begin
        if (reset) begin
            cnt       <= 3'd0;
            pulse_cnt <= 2'd0;
            out       <= 1'b0;
            fired     <= 1'b0;
        end else begin
            if (fired) begin
                // �Ѿ���������ϵͳ������ֱ�� reset
                out <= 1'b0;
            end else begin
                if (out) begin
                    // out �Ѿ�Ϊ 1������������
                    if (pulse_cnt == 2'd1) begin
                        out       <= 1'b0;
                        fired     <= 1'b1;
                        pulse_cnt <= 2'd0;
                    end else begin
                        pulse_cnt <= pulse_cnt + 2'd1;
                        out       <= 1'b1;
                    end
                end else begin
                    // out == 0����δ����
                    if (in && data) begin
                        if (cnt == 3'd3) begin
                            out       <= 1'b1;   // ���� 4 clk �󴥷�
                            pulse_cnt <= 2'd0;
                            cnt       <= cnt;    // ����
                        end else begin
                            cnt <= cnt + 3'd1;
                        end
                    end else begin
                        cnt <= 3'd0;  // ��һΪ 0�����¼���
                    end
                end
            end
        end
    end

endmodule
