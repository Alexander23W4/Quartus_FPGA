library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- �޸�ʵ������������֮ǰ��multiplier_4x4��ͻ
entity bcd_multiplier is
    port(
        a, b : in  std_logic_vector(3 downto 0);  -- 4λ����
        bcd_hundreds : out std_logic_vector(3 downto 0);  -- ��λBCD (0-2)
        bcd_tens     : out std_logic_vector(3 downto 0);  -- ʮλBCD (0-9)
        bcd_ones     : out std_logic_vector(3 downto 0)   -- ��λBCD (0-9)
    );
end entity;

architecture behavioral of bcd_multiplier is
    signal product : unsigned(7 downto 0);  -- ԭʼ�˻�
begin
    -- ����˻�
    product <= unsigned(a) * unsigned(b);
    
    -- ������תBCD
    process(product)
        variable bcd_temp : unsigned(11 downto 0);  -- 3��BCD�빲12λ
    begin
        -- ��ʼ��
        bcd_temp := (others => '0');
        bcd_temp(7 downto 0) := product;
        
        -- ˫����ת����8��ѭ����
        for i in 0 to 7 loop
            -- ��λ����
            if bcd_temp(11 downto 8) >= 5 then
                bcd_temp(11 downto 8) := bcd_temp(11 downto 8) + 3;
            end if;
            
            -- ʮλ����
            if bcd_temp(7 downto 4) >= 5 then
                bcd_temp(7 downto 4) := bcd_temp(7 downto 4) + 3;
            end if;
            
            -- ��λ����
            if bcd_temp(3 downto 0) >= 5 then
                bcd_temp(3 downto 0) := bcd_temp(3 downto 0) + 3;
            end if;
            
            -- ����
            bcd_temp := bcd_temp(10 downto 0) & '0';
        end loop;
        
        -- ���BCD��
        bcd_hundreds <= std_logic_vector(bcd_temp(11 downto 8));  -- ��λ
        bcd_tens     <= std_logic_vector(bcd_temp(7 downto 4));   -- ʮλ
        bcd_ones     <= std_logic_vector(bcd_temp(3 downto 0));   -- ��λ
    end process;
end architecture;

-- �򻯰棨�������㣬��ֱ�ۣ�
architecture simple of bcd_multiplier is
    signal product_int : integer range 0 to 255;
begin
    -- ����˻�
    product_int <= to_integer(unsigned(a)) * to_integer(unsigned(b));
    
    -- ֱ�Ӽ����λ��ʮλ����λ
    process(product_int)
        variable hundreds, tens, ones : integer range 0 to 9;
    begin
        -- �����λ����
        hundreds := product_int / 100;
        tens     := (product_int / 10) mod 10;
        ones     := product_int mod 10;
        
        -- ת��Ϊ������
        bcd_hundreds <= std_logic_vector(to_unsigned(hundreds, 4));
        bcd_tens     <= std_logic_vector(to_unsigned(tens, 4));
        bcd_ones     <= std_logic_vector(to_unsigned(ones, 4));
    end process;
end architecture;