library ieee;
use ieee.std_logic_1164.all;

-- 4λ�����Ĵ���������ȫ���ֿ���
entity latch_4bit_separate is
    port (
        -- ʱ�Ӻ�ʹ��
        clk      : in std_logic;        -- ʱ�ӣ�����ʱ��ʱ�ɽӸߵ�ƽ��
        set      : in std_logic;        -- ��λʹ�ܣ�����Ч��
        clear    : in std_logic;        -- ���㣨����Ч��
        
        -- 4λ���루�ֿ������ţ�
        din0     : in std_logic;        -- ����λ0
        din1     : in std_logic;        -- ����λ1  
        din2     : in std_logic;        -- ����λ2
        din3     : in std_logic;        -- ����λ3
        
        -- 4λ������ֿ������ţ�
        dout0    : out std_logic;       -- ���λ0
        dout1    : out std_logic;       -- ���λ1
        dout2    : out std_logic;       -- ���λ2
        dout3    : out std_logic        -- ���λ3
    );
end entity latch_4bit_separate;

architecture behavioral of latch_4bit_separate is
    -- �ڲ��Ĵ���λ
    signal reg0, reg1, reg2, reg3 : std_logic := '0';
    
    -- �����ź�
    signal fb0, fb1, fb2, fb3 : std_logic;
begin
    -- �����߼���������������ֵ
    fb0 <= din0 or reg0;
    fb1 <= din1 or reg1;
    fb2 <= din2 or reg2;
    fb3 <= din3 or reg3;
    
    -- 4��������D���������൱��4��7474��
    -- λ0������
    process(clk, clear)
    begin
        if clear = '1' then
            reg0 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg0 <= fb0;
            end if;
        end if;
    end process;
    
    -- λ1������
    process(clk, clear)
    begin
        if clear = '1' then
            reg1 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg1 <= fb1;
            end if;
        end if;
    end process;
    
    -- λ2������
    process(clk, clear)
    begin
        if clear = '1' then
            reg2 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg2 <= fb2;
            end if;
        end if;
    end process;
    
    -- λ3������
    process(clk, clear)
    begin
        if clear = '1' then
            reg3 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg3 <= fb3;
            end if;
        end if;
    end process;
    
    -- �������
    dout0 <= reg0;
    dout1 <= reg1;
    dout2 <= reg2;
    dout3 <= reg3;
end architecture behavioral;

-- ���򵥵ĵ�ƽ�����汾������Ҫʱ�ӣ�
architecture simple of latch_4bit_separate is
    signal q0, q1, q2, q3 : std_logic := '0';
begin
    -- λ0��һ������Ϊ1�����棬ֱ������
    process(set, clear, din0)
    begin
        if clear = '1' then
            q0 <= '0';
        elsif set = '1' and din0 = '1' then
            q0 <= '1';
        end if;
    end process;
    
    -- λ1
    process(set, clear, din1)
    begin
        if clear = '1' then
            q1 <= '0';
        elsif set = '1' and din1 = '1' then
            q1 <= '1';
        end if;
    end process;
    
    -- λ2
    process(set, clear, din2)
    begin
        if clear = '1' then
            q2 <= '0';
        elsif set = '1' and din2 = '1' then
            q2 <= '1';
        end if;
    end process;
    
    -- λ3
    process(set, clear, din3)
    begin
        if clear = '1' then
            q3 <= '0';
        elsif set = '1' and din3 = '1' then
            q3 <= '1';
        end if;
    end process;
    
    -- ���
    dout0 <= q0;
    dout1 <= q1;
    dout2 <= q2;
    dout3 <= q3;
end architecture simple;

-- ʹ��ʾ��
architecture usage_example of latch_4bit_separate is
begin
    -- ��򵥵��÷���clk�Ӹߵ�ƽ��set����
    -- ����ֻҪ������Ϊ1����������
end architecture usage_example;