library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bcd_mult4x4 is
    port(
        a, b : in  std_logic_vector(3 downto 0);  -- 4λ����
        bcd2 : out std_logic_vector(3 downto 0);  -- ��λBCD (0-2)
        bcd1 : out std_logic_vector(3 downto 0);  -- ʮλBCD (0-9)
        bcd0 : out std_logic_vector(3 downto 0)   -- ��λBCD (0-9)
    );
end entity;

architecture behavioral of bcd_mult4x4 is
    signal product : unsigned(7 downto 0);  -- ԭʼ�˻�
    signal temp    : unsigned(7 downto 0);  -- ת������ʱ����
begin
    -- ����˻�
    product <= unsigned(a) * unsigned(b);
    
    -- ������תBCD (˫����)
    process(product)
        variable bcd_temp : unsigned(11 downto 0);  -- 3��BCD�빲12λ
    begin
        -- ��ʼ��
        bcd_temp := (others => '0');
        bcd_temp(7 downto 0) := product;
        
        -- ѭ��8�Σ�ÿ����λ������BCD
        for i in 0 to 7 loop
            -- ����λ�Ƿ�>=5
            if bcd_temp(11 downto 8) >= 5 then
                bcd_temp(11 downto 8) := bcd_temp(11 downto 8) + 3;
            end if;
            
            -- ���ʮλ�Ƿ�>=5
            if bcd_temp(7 downto 4) >= 5 then
                bcd_temp(7 downto 4) := bcd_temp(7 downto 4) + 3;
            end if;
            
            -- ����λ�Ƿ�>=5
            if bcd_temp(3 downto 0) >= 5 then
                bcd_temp(3 downto 0) := bcd_temp(3 downto 0) + 3;
            end if;
            
            -- ����һλ
            bcd_temp := bcd_temp(10 downto 0) & '0';
        end loop;
        
        -- ���BCD��
        bcd2 <= std_logic_vector(bcd_temp(11 downto 8));  -- ��λ
        bcd1 <= std_logic_vector(bcd_temp(7 downto 4));   -- ʮλ
        bcd0 <= std_logic_vector(bcd_temp(3 downto 0));   -- ��λ
    end process;
end architecture;

-- �򻯰棨�����Χֻ��0-99������Ҫ��λ����
architecture simple of bcd_mult4x4 is
    signal product : integer range 0 to 255;
begin
    product <= to_integer(unsigned(a)) * to_integer(unsigned(b));
    
    bcd2 <= "0000" when product < 100 else  -- ��λ����0��1
            "0001" when product < 200 else
            "0010";
    
    bcd1 <= std_logic_vector(to_unsigned((product / 10) mod 10, 4));
    bcd0 <= std_logic_vector(to_unsigned(product mod 10, 4));
end architecture;