library ieee;
use ieee.std_logic_1164.all;

-- 8λ�����Ĵ���������ȫ���ֿ���
entity latch_8bit_separate is
    port (
        -- ʱ�Ӻ�ʹ��
        clk      : in std_logic;        -- ʱ�ӣ�����ʱ��ʱ�ɽӸߵ�ƽ��
        set      : in std_logic;        -- ��λʹ�ܣ�����Ч��
        clear    : in std_logic;        -- ���㣨����Ч��
        
        -- 8λ���루�ֿ������ţ�
        din0     : in std_logic;        -- ����λ0
        din1     : in std_logic;        -- ����λ1  
        din2     : in std_logic;        -- ����λ2
        din3     : in std_logic;        -- ����λ3
        din4     : in std_logic;        -- ����λ4
        din5     : in std_logic;        -- ����λ5
        din6     : in std_logic;        -- ����λ6
        din7     : in std_logic;        -- ����λ7
        
        -- 8λ������ֿ������ţ�
        dout0    : out std_logic;       -- ���λ0
        dout1    : out std_logic;       -- ���λ1
        dout2    : out std_logic;       -- ���λ2
        dout3    : out std_logic;       -- ���λ3
        dout4    : out std_logic;       -- ���λ4
        dout5    : out std_logic;       -- ���λ5
        dout6    : out std_logic;       -- ���λ6
        dout7    : out std_logic        -- ���λ7
    );
end entity latch_8bit_separate;

architecture behavioral of latch_8bit_separate is
    -- �ڲ��Ĵ���λ
    signal reg0, reg1, reg2, reg3, reg4, reg5, reg6, reg7 : std_logic := '0';
    
    -- �����ź�
    signal fb0, fb1, fb2, fb3, fb4, fb5, fb6, fb7 : std_logic;
begin
    -- �����߼���������������ֵ
    fb0 <= din0 or reg0;
    fb1 <= din1 or reg1;
    fb2 <= din2 or reg2;
    fb3 <= din3 or reg3;
    fb4 <= din4 or reg4;
    fb5 <= din5 or reg5;
    fb6 <= din6 or reg6;
    fb7 <= din7 or reg7;
    
    -- 8��������D���������൱��8��7474��
    
    -- λ0������
    process(clk, clear)
    begin
        if clear = '1' then
            reg0 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg0 <= fb0;
            end if;
        end if;
    end process;
    
    -- λ1������
    process(clk, clear)
    begin
        if clear = '1' then
            reg1 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg1 <= fb1;
            end if;
        end if;
    end process;
    
    -- λ2������
    process(clk, clear)
    begin
        if clear = '1' then
            reg2 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg2 <= fb2;
            end if;
        end if;
    end process;
    
    -- λ3������
    process(clk, clear)
    begin
        if clear = '1' then
            reg3 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg3 <= fb3;
            end if;
        end if;
    end process;
    
    -- λ4������
    process(clk, clear)
    begin
        if clear = '1' then
            reg4 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg4 <= fb4;
            end if;
        end if;
    end process;
    
    -- λ5������
    process(clk, clear)
    begin
        if clear = '1' then
            reg5 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg5 <= fb5;
            end if;
        end if;
    end process;
    
    -- λ6������
    process(clk, clear)
    begin
        if clear = '1' then
            reg6 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg6 <= fb6;
            end if;
        end if;
    end process;
    
    -- λ7������
    process(clk, clear)
    begin
        if clear = '1' then
            reg7 <= '0';
        elsif rising_edge(clk) then
            if set = '1' then
                reg7 <= fb7;
            end if;
        end if;
    end process;
    
    -- �������
    dout0 <= reg0;
    dout1 <= reg1;
    dout2 <= reg2;
    dout3 <= reg3;
    dout4 <= reg4;
    dout5 <= reg5;
    dout6 <= reg6;
    dout7 <= reg7;
end architecture behavioral;

-- ���򵥵ĵ�ƽ�����汾���Ƽ���
architecture simple of latch_8bit_separate is
    signal q0, q1, q2, q3, q4, q5, q6, q7 : std_logic := '0';
begin
    -- λ0��һ������Ϊ1�����棬ֱ������
    process(set, clear, din0)
    begin
        if clear = '1' then
            q0 <= '0';
        elsif set = '1' and din0 = '1' then
            q0 <= '1';
        end if;
    end process;
    
    -- λ1
    process(set, clear, din1)
    begin
        if clear = '1' then
            q1 <= '0';
        elsif set = '1' and din1 = '1' then
            q1 <= '1';
        end if;
    end process;
    
    -- λ2
    process(set, clear, din2)
    begin
        if clear = '1' then
            q2 <= '0';
        elsif set = '1' and din2 = '1' then
            q2 <= '1';
        end if;
    end process;
    
    -- λ3
    process(set, clear, din3)
    begin
        if clear = '1' then
            q3 <= '0';
        elsif set = '1' and din3 = '1' then
            q3 <= '1';
        end if;
    end process;
    
    -- λ4
    process(set, clear, din4)
    begin
        if clear = '1' then
            q4 <= '0';
        elsif set = '1' and din4 = '1' then
            q4 <= '1';
        end if;
    end process;
    
    -- λ5
    process(set, clear, din5)
    begin
        if clear = '1' then
            q5 <= '0';
        elsif set = '1' and din5 = '1' then
            q5 <= '1';
        end if;
    end process;
    
    -- λ6
    process(set, clear, din6)
    begin
        if clear = '1' then
            q6 <= '0';
        elsif set = '1' and din6 = '1' then
            q6 <= '1';
        end if;
    end process;
    
    -- λ7
    process(set, clear, din7)
    begin
        if clear = '1' then
            q7 <= '0';
        elsif set = '1' and din7 = '1' then
            q7 <= '1';
        end if;
    end process;
    
    -- ���
    dout0 <= q0;
    dout1 <= q1;
    dout2 <= q2;
    dout3 <= q3;
    dout4 <= q4;
    dout5 <= q5;
    dout6 <= q6;
    dout7 <= q7;
end architecture simple;

-- �򻯰汾2��ʹ��generate���
architecture compact of latch_8bit_separate is
    type reg_array is array (0 to 7) of std_logic;
    signal q : reg_array := (others => '0');
	signal d : reg_array;  -- ��Ϊ���
begin
    -- ��������
    d(0) <= din0;
    d(1) <= din1;
    d(2) <= din2;
    d(3) <= din3;
    d(4) <= din4;
    d(5) <= din5;
    d(6) <= din6;
    d(7) <= din7;
    
    -- ����8��������
    gen_latch: for i in 0 to 7 generate
        process(set, clear, d(i))
        begin
            if clear = '1' then
                q(i) <= '0';
            elsif set = '1' and d(i) = '1' then
                q(i) <= '1';
            end if;
        end process;
    end generate;
    
    -- ���
    dout0 <= q(0);
    dout1 <= q(1);
    dout2 <= q(2);
    dout3 <= q(3);
    dout4 <= q(4);
    dout5 <= q(5);
    dout6 <= q(6);
    dout7 <= q(7);
end architecture compact;